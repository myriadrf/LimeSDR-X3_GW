-- ----------------------------------------------------------------------------	
-- FILE:	cdcmcfg.vhd
-- DESCRIPTION:	Serial configuration interface to control TX modules
-- DATE:	March 16, 2021
-- AUTHOR(s):	Lime Microsystems
-- REVISIONS:	
-- ----------------------------------------------------------------------------	

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mem_package.all;
use work.revisions.all;
use work.cdcmcfg_pkg.all;

-- ----------------------------------------------------------------------------
-- Entity declaration
-- ----------------------------------------------------------------------------
entity cdcmcfg is
   generic (
   CDCM_REG_0_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_1_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_2_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_3_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_4_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_5_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_6_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_7_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_8_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_9_DEFAULT  : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_10_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_11_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_12_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_13_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_14_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_15_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_16_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_17_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_18_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_19_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000";
   CDCM_REG_20_DEFAULT : std_logic_vector(15 downto 0) := B"0000_0000_0000_0000"
   );
   port (
      -- Address and location of this module
      -- Will be hard wired at the top level
      maddress    : in  std_logic_vector(9 downto 0);
      mimo_en     : in  std_logic;   -- MIMO enable, from TOP SPI (always 1)
   
      -- Serial port IOs
      sdin        : in  std_logic;  -- Data in
      sclk        : in  std_logic;  -- Data clock
      sen         : in  std_logic;  -- Enable signal (active low)
      sdout       : out std_logic;  -- Data out
   
      -- Signals coming from the pins or top level serial interface
      lreset      : in  std_logic;  -- Logic reset signal, resets logic cells only  (use only one reset)
      mreset      : in  std_logic;  -- Memory reset signal, resets configuration memory only (use only one reset)
      
      oen         : out std_logic;  --nc
      stateo      : out std_logic_vector(5 downto 0)
--      stateo      : out std_logic_vector(5 downto 0);
--      to_cdcmcfg  : in  t_TO_CDCMCFG;
--      from_cdcmcfg: out t_FROM_CDCMCFG
      
      
   );
end cdcmcfg;

-- ----------------------------------------------------------------------------
-- Architecture
-- ----------------------------------------------------------------------------
architecture cdcmcfg_arch of cdcmcfg is

   signal inst_reg: std_logic_vector(15 downto 0);    -- Instruction register
   signal inst_reg_en: std_logic;

   signal din_reg: std_logic_vector(15 downto 0);     -- Data in register
   signal din_reg_en: std_logic;
   
   signal dout_reg: std_logic_vector(15 downto 0);    -- Data out register
   signal dout_reg_sen, dout_reg_len: std_logic;
   
   signal mem: marray32x16;                           -- Config memory
   signal mem_we: std_logic;
   
   signal oe: std_logic;                              -- Tri state buffers control
   signal spi_config_data_rev	: std_logic_vector(143 downto 0);
      
   -- Components
   use work.mcfg_components.mcfg32wm_fsm;
   for all: mcfg32wm_fsm use entity work.mcfg32wm_fsm(mcfg32wm_fsm_arch);

begin

   -- ---------------------------------------------------------------------------------------------
   -- Finite state machines
   -- ---------------------------------------------------------------------------------------------
   fsm: mcfg32wm_fsm port map( 
      address => maddress, mimo_en => mimo_en, inst_reg => inst_reg, sclk => sclk, sen => sen, reset => lreset,
      inst_reg_en => inst_reg_en, din_reg_en => din_reg_en, dout_reg_sen => dout_reg_sen,
      dout_reg_len => dout_reg_len, mem_we => mem_we, oe => oe, stateo => stateo);
      
   -- ---------------------------------------------------------------------------------------------
   -- Instruction register
   -- ---------------------------------------------------------------------------------------------
   inst_reg_proc: process(sclk, lreset)
      variable i: integer;
   begin
      if lreset = '0' then
         inst_reg <= (others => '0');
      elsif sclk'event and sclk = '1' then
         if inst_reg_en = '1' then
            for i in 15 downto 1 loop
               inst_reg(i) <= inst_reg(i-1);
            end loop;
            inst_reg(0) <= sdin;
         end if;
      end if;
   end process inst_reg_proc;

   -- ---------------------------------------------------------------------------------------------
   -- Data input register
   -- ---------------------------------------------------------------------------------------------
   din_reg_proc: process(sclk, lreset)
      variable i: integer;
   begin
      if lreset = '0' then
         din_reg <= (others => '0');
      elsif sclk'event and sclk = '1' then
         if din_reg_en = '1' then
            for i in 15 downto 1 loop
               din_reg(i) <= din_reg(i-1);
            end loop;
            din_reg(0) <= sdin;
         end if;
      end if;
   end process din_reg_proc;

   -- ---------------------------------------------------------------------------------------------
   -- Data output register
   -- ---------------------------------------------------------------------------------------------
   dout_reg_proc: process(sclk, lreset)
      variable i: integer;
   begin
      if lreset = '0' then
         dout_reg <= (others => '0');
      elsif sclk'event and sclk = '0' then
         -- Shift operation
         if dout_reg_sen = '1' then
            for i in 15 downto 1 loop
               dout_reg(i) <= dout_reg(i-1);
            end loop;
            dout_reg(0) <= dout_reg(15);
         -- Load operation
         elsif dout_reg_len = '1' then
            case inst_reg(4 downto 0) is  -- mux read-only outputs
               when others  => dout_reg <= mem(to_integer(unsigned(inst_reg(4 downto 0))));
            end case;
         end if;
      end if;
   end process dout_reg_proc;
   
   -- Tri state buffer to connect multiple serial interfaces in parallel
   --sdout <= dout_reg(7) when oe = '1' else 'Z';

-- sdout <= dout_reg(7);
-- oen <= oe;

   sdout <= dout_reg(15) and oe;
   oen <= oe;
   -- ---------------------------------------------------------------------------------------------
   -- Configuration memory
   -- --------------------------------------------------------------------------------------------- 
   ram: process(sclk, mreset) --(remap)
   begin
      -- Defaults
      if mreset = '0' then
         mem(0)   <= CDCM_REG_0_DEFAULT ;  -- 00 free, CDCM_REG_0
         mem(1)   <= CDCM_REG_1_DEFAULT ;  -- 00 free, CDCM_REG_1
         mem(2)   <= CDCM_REG_2_DEFAULT ;  -- 00 free, CDCM_REG_2
         mem(3)   <= CDCM_REG_3_DEFAULT ;  -- 00 free, CDCM_REG_3
         mem(4)   <= CDCM_REG_4_DEFAULT ;  -- 00 free, CDCM_REG_4
         mem(5)   <= CDCM_REG_5_DEFAULT ;  -- 00 free, CDCM_REG_5
         mem(6)   <= CDCM_REG_6_DEFAULT ;  -- 00 free, CDCM_REG_6
         mem(7)   <= CDCM_REG_7_DEFAULT ;  -- 00 free, CDCM_REG_7
         mem(8)   <= CDCM_REG_8_DEFAULT ;  -- 00 free, CDCM_REG_8
         mem(9)   <= CDCM_REG_9_DEFAULT ;  -- 00 free, CDCM_REG_9
         mem(10)  <= CDCM_REG_10_DEFAULT;  -- 00 free, CDCM_REG_10
         mem(11)  <= CDCM_REG_11_DEFAULT;  -- 00 free, CDCM_REG_11
         mem(12)  <= CDCM_REG_12_DEFAULT;  -- 00 free, CDCM_REG_12
         mem(13)  <= CDCM_REG_13_DEFAULT;  -- 00 free, CDCM_REG_13
         mem(14)  <= CDCM_REG_14_DEFAULT;  -- 00 free, CDCM_REG_14
         mem(15)  <= CDCM_REG_15_DEFAULT;  -- 00 free, CDCM_REG_15
         mem(16)  <= CDCM_REG_16_DEFAULT;  -- 00 free, CDCM_REG_16
         mem(17)  <= CDCM_REG_17_DEFAULT;  -- 00 free, CDCM_REG_17
         mem(18)  <= CDCM_REG_18_DEFAULT;  -- 00 free, CDCM_REG_18
         mem(19)  <= CDCM_REG_19_DEFAULT;  -- 00 free, CDCM_REG_19
         mem(20)  <= CDCM_REG_20_DEFAULT;  -- 00 free, CDCM_REG_20
         mem(21)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED(15:3), CDCM_CONFIG_ERROR ,CDCM_CONFIG_DONE, CDCM_CONFIG_START
         mem(22)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(23)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(24)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(25)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(26)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(27)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(28)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(29)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(30)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         mem(31)  <= "0000000000000000";  -- 00 free, UNUSED/RESERVED
         
      elsif sclk'event and sclk = '1' then
            if mem_we = '1' then
               mem(to_integer(unsigned(inst_reg(4 downto 0)))) <= din_reg(14 downto 0) & sdin;
            end if;
            
            if dout_reg_len = '0' then
--               for_loop : for i in 0 to 3 loop
--                  mem(3)(i+4) <= not mem(3)(i);
--               end loop;
            end if;
            
      end if;
   end process ram;
   
   -- ---------------------------------------------------------------------------------------------
   -- Decoding logic
   -- ---------------------------------------------------------------------------------------------

--empty


end cdcmcfg_arch;
